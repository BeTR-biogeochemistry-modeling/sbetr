netcdf uniform_steadystate_grid {
dimensions:
	levgrnd = 15 ;
	lndgrid = 1 ;
variables:
	double BSW(levgrnd, lndgrid) ;
		BSW:long_name = "slope of soil water retention curve" ;
		BSW:units = "unitless" ;
		BSW:_FillValue = 9.9999996169031625e+35 ;
		BSW:missing_value = 9.99999962e+35f ;
	double DZSOI(levgrnd, lndgrid) ;
		DZSOI:long_name = "soil thickness" ;
		DZSOI:units = "m" ;
		DZSOI:_FillValue = 9.9999996169031625e+35 ;
		DZSOI:missing_value = 9.99999962e+35f ;
	double WATSAT(levgrnd, lndgrid) ;
		WATSAT:long_name = "saturated soil water content (porosity)" ;
		WATSAT:units = "mm3/mm3" ;
		WATSAT:_FillValue = 9.9999996169031625e+35 ;
		WATSAT:missing_value = 9.99999962e+35f ;
	double ZSOI(levgrnd, lndgrid) ;
		ZSOI:long_name = "soil depth" ;
		ZSOI:units = "m" ;
		ZSOI:_FillValue = 9.9999996169031625e+35 ;
		ZSOI:missing_value = 9.99999962e+35f ;
	double lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 9.9999996169031625e+35 ;
		lat:missing_value = 9.99999962e+35f ;
	double levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	double lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 9.9999996169031625e+35 ;
		lon:missing_value = 9.99999962e+35f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "Tue Jan 26 14:08:50 2016: ncks -v WATSAT,lon,lat,DZSOI,ZSOI,BSW CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15.clm2.h0.0001-01-01-00000.nc sierra_grid.nc\n",
			"created on 01/20/16 13:41:24" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "lawrencium-lr3" ;
		:username = "jitang" ;
		:version = "cesm1_3_beta10" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15" ;
		:Surface_dataset = "surfdata_US-Blo_grid_c160115.nc" ;
		:Initial_conditions_dataset = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.2016-01-15.clm2.r.0061-01-01-00000.nc" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:NCO = "\"4.5.3\"" ;
data:

 BSW =
  5.5819539999999996,
  5.8422970000000003,
  6.1484259999999997,
  6.3773369999999998,
  6.7252010000000002,
  6.8982460000000003,
  7.3739509999999999,
  7.2094379999999996,
  7.2030000000000003,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996 ;

 DZSOI =
  0.017512819999999998,
  0.027578970000000001,
  0.045470030000000002,
  0.074967409999999998,
  0.1236004,
  0.20378260000000001,
  0.33598060000000002,
  0.55393840000000005,
  0.91329000000000005,
  1.5057609999999999,
  2.48258,
  4.0930819999999999,
  6.7483510000000004,
  11.126150000000001,
  13.851150000000001 ;

 WATSAT =
  0.50330949999999997,
  0.46785690000000002,
  0.44546940000000002,
  0.4358359,
  0.43314900000000001,
  0.42817480000000002,
  0.42955460000000001,
  0.42528389999999999,
  0.42348000000000002,
  0.42852000000000001,
  0.42852000000000001,
  0.42852000000000001,
  0.42852000000000001,
  0.42852000000000001,
  0.42852000000000001 ;

 ZSOI =
  0.0071006350000000001,
  0.027924999999999998,
  0.062258580000000001,
  0.1188651,
  0.2121934,
  0.3660658,
  0.61975849999999999,
  1.038027,
  1.727635,
  2.8646069999999999,
  4.7391569999999996,
  7.8297660000000002,
  12.925319999999999,
  21.32647,
  35.177619999999997 ;

 lat = 38.895200000000003 ;

 levgrnd = 0.0071006350000000001, 0.027924999999999998, 0.062258580000000001, 
    0.1188651, 0.2121934, 0.3660658, 0.61975849999999999, 1.038027, 1.727635, 
    2.8646069999999999, 4.7391569999999996, 7.8297660000000002, 
    12.925319999999999, 21.32647, 35.177619999999997 ;

 lon = 239.3673 ;
}
