netcdf uniform_steadystate_grid {
dimensions:
	levgrnd = 15 ;
	lndgrid = 1 ;
variables:
	float BSW(levgrnd, lndgrid) ;
		BSW:long_name = "slope of soil water retention curve" ;
		BSW:units = "unitless" ;
		BSW:_FillValue = 1.e+36f ;
		BSW:missing_value = 1.e+36f ;
	float DZSOI(levgrnd, lndgrid) ;
		DZSOI:long_name = "soil thickness" ;
		DZSOI:units = "m" ;
		DZSOI:_FillValue = 1.e+36f ;
		DZSOI:missing_value = 1.e+36f ;
	float WATSAT(levgrnd, lndgrid) ;
		WATSAT:long_name = "saturated soil water content (porosity)" ;
		WATSAT:units = "mm3/mm3" ;
		WATSAT:_FillValue = 1.e+36f ;
		WATSAT:missing_value = 1.e+36f ;
	float ZSOI(levgrnd, lndgrid) ;
		ZSOI:long_name = "soil depth" ;
		ZSOI:units = "m" ;
		ZSOI:_FillValue = 1.e+36f ;
		ZSOI:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "Tue Jan 26 14:08:50 2016: ncks -v WATSAT,lon,lat,DZSOI,ZSOI,BSW CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15.clm2.h0.0001-01-01-00000.nc sierra_grid.nc\n",
			"created on 01/20/16 13:41:24" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "lawrencium-lr3" ;
		:username = "jitang" ;
		:version = "cesm1_3_beta10" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.norm.2016-01-15" ;
		:Surface_dataset = "surfdata_US-Blo_grid_c160115.nc" ;
		:Initial_conditions_dataset = "CLM_USRDAT.ICLM45.lawrencium-lr3.intel.5656685.2016-01-15.clm2.r.0061-01-01-00000.nc" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:NCO = "\"4.5.3\"" ;
data:

 BSW =
  5.581954,
  5.842297,
  6.148426,
  6.377337,
  6.725201,
  6.898246,
  7.373951,
  7.209438,
  7.203,
  8.475,
  8.475,
  8.475,
  8.475,
  8.475,
  8.475 ;

 DZSOI =
  0.01751282,
  0.02757897,
  0.04547003,
  0.07496741,
  0.1236004,
  0.2037826,
  0.3359806,
  0.5539384,
  0.91329,
  1.505761,
  2.48258,
  4.093082,
  6.748351,
  11.12615,
  13.85115 ;

 WATSAT =
  0.5033095,
  0.4678569,
  0.4454694,
  0.4358359,
  0.433149,
  0.4281748,
  0.4295546,
  0.4252839,
  0.42348,
  0.42852,
  0.42852,
  0.42852,
  0.42852,
  0.42852,
  0.42852 ;

 ZSOI =
  0.007100635,
  0.027925,
  0.06225858,
  0.1188651,
  0.2121934,
  0.3660658,
  0.6197585,
  1.038027,
  1.727635,
  2.864607,
  4.739157,
  7.829766,
  12.92532,
  21.32647,
  35.17762 ;

 lat = 38.8952 ;

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 lon = 239.3673 ;
}
