netcdf sierra_steadystate {
dimensions:
	levgrnd = 15 ;
	lndgrid = 1 ;
	time = 1 ;
variables:
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:units = "K" ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:missing_value = 1.e+36f ;
		TSOI:_FillValue = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:missing_value = 1.e+36f ;
		H2OSOI:_FillValue = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:units = "kg/m2" ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:missing_value = 1.e+36f ;
		SOILICE:_FillValue = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:units = "Pa" ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:missing_value = 1.e+36f ;
		PBOT:_FillValue = 1.e+36f ;
	float QFLX_ROOTSOI(time, levgrnd, lndgrid) ;
		QFLX_ROOTSOI:units = "m/s" ;
		QFLX_ROOTSOI:long_name = "depth dependent root water uptake" ;
		QFLX_ROOTSOI:cell_methods = "time: mean" ;
		QFLX_ROOTSOI:missing_value = 1.e+36f ;
		QFLX_ROOTSOI:_FillValue = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:units = "K" ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:missing_value = 1.e+36f ;
		TBOT:_FillValue = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:missing_value = 1.e+36f ;
		QCHARGE:_FillValue = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:units = "mm/s" ;
		QINFL:long_name = "infiltration" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:missing_value = 1.e+36f ;
		QINFL:_FillValue = 1.e+36f ;
	float time(time) ;
                time:long_name = "time" ;
                time:units = "days since 0001-01-01 00:00:00" ;
                time:calendar = "noleap" ;
                time:bounds = "time_bounds" ;
data:

 TSOI =
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0,
  283.0 ;

 H2OSOI =
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3,
  0.3 ;

 SOILICE =
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0,
  0 ;

 QFLX_ROOTSOI =
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10,
  3.0e-10 ;

 PBOT =
  101325.0 ;

 TBOT =
  278.0 ;

 QCHARGE =
  1.0e-05 ;

 QINFL =
  4.0e-05 ;

 time = 1.0 ;
}
