netcdf uniform_steadystate_grid.cdl {
dimensions:
	levgrnd = 15 ;
	lndgrid = 1 ;
variables:
	double BSW(levgrnd, lndgrid) ;
		BSW:long_name = "slope of soil water retention curve" ;
		BSW:units = "unitless" ;
		BSW:_FillValue = 9.9999996169031625e+35 ;
		BSW:missing_value = 9.99999962e+35f ;
	double WATSAT(levgrnd, lndgrid) ;
		WATSAT:long_name = "saturated soil water content (porosity)" ;
		WATSAT:units = "mm3/mm3" ;
		WATSAT:_FillValue = 9.9999996169031625e+35 ;
		WATSAT:missing_value = 9.99999962e+35f ;

// global attributes:
		:title = "Standalone BeTR uniform soil parameters." ;
		:comment = "NOTE(bja, 201604) created by arbitrarily removing variability from another file!" ;
		:Conventions = "CF-1.0" ;
data:

 BSW =
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996,
  8.4749999999999996 ;

 WATSAT =
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5,
  0.5 ;
}
